module Wire(
input logic a, output logic z
    );
    assign z=a;
endmodule
